
module top (a, b, y);
input y;
output a, b;

buf(a, b, y);

endmodule
