

module top (a, b, y);
input y;
output a, b;

not(a, b, y);

endmodule
